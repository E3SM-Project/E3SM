netcdf clm_exp_grid.cdl {
dimensions:
	levgrnd = 15 ;
	lndgrid = 1 ;
variables:
	double BSW(levgrnd, lndgrid) ;
		BSW:long_name = "slope of soil water retention curve" ;
		BSW:units = "unitless" ;
		BSW:_FillValue = 9.99999961690316e+35 ;
		BSW:missing_value = 1.e+36f ;
	double SUCSAT(levgrnd, lndgrid) ;
		SUCSAT:long_name = "saturated soil matric potential" ;
		SUCSAT:units = "mm" ;
		SUCSAT:_FillValue = 1.e+36f ;
		SUCSAT:missing_value = 1.e+36f ;
	double DZSOI(levgrnd, lndgrid) ;
		DZSOI:long_name = "soil thickness" ;
		DZSOI:units = "m" ;
		DZSOI:_FillValue = 9.99999961690316e+35 ;
		DZSOI:missing_value = 1.e+36f ;
	double PCTSAND(levgrnd, lndgrid) ;
		PCTSAND:long_name = "percentage of sand" ;
		PCTSAND:units = "%" ;
		PCTSAND:_FillValue = 9.99999961690316e+35 ;
		PCTSAND:missing_value = 1.e+36f ;
	double WATSAT(levgrnd, lndgrid) ;
		WATSAT:long_name = "saturated soil water content (porosity)" ;
		WATSAT:units = "mm3/mm3" ;
		WATSAT:_FillValue = 9.99999961690316e+35 ;
		WATSAT:missing_value = 1.e+36f ;
	double ZSOI(levgrnd, lndgrid) ;
		ZSOI:long_name = "soil depth" ;
		ZSOI:units = "m" ;
		ZSOI:_FillValue = 9.99999961690316e+35 ;
		ZSOI:missing_value = 1.e+36f ;
	double lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 9.99999961690316e+35 ;
		lat:missing_value = 1.e+36f ;
	double levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	double lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 9.99999961690316e+35 ;
		lon:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "Tue Jan 26 14:08:50 2016: ncks -v WATSAT,lon,lat,DZSOI,ZSOI,BSW CLM_USRDAT.ICLM45.lawrencium-lr3.intel.5656685.norm.2016-01-15.clm2.h0.0001-01-01-00000.nc sierra_grid.nc\n",
			"created on 01/20/16 13:41:24" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "lawrencium-lr3" ;
		:username = "jitang" ;
		:version = "cesm1_3_beta10" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "CLM_USRDAT.ICLM45.lawrencium-lr3.intel.5656685.norm.2016-01-15" ;
		:Surface_dataset = "surfdata_US-Blo_grid_c160115.nc" ;
		:Initial_conditions_dataset = "CLM_USRDAT.ICLM45.lawrencium-lr3.intel.5656685.2016-01-15.clm2.r.0061-01-01-00000.nc" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:NCO = "\"4.5.3\"" ;
data:

 BSW =
  5.581954,
  5.8422966,
  6.14842558,
  6.3773365,
  6.72520113,
  6.89824629,
  7.37395144,
  7.20943785,
  7.20300007,
  8.47500038,
  8.47500038,
  8.47500038,
  8.47500038,
  8.47500038,
  8.47500038 ;

 SUCSAT =
  139.0655,
  149.7077,
  156.4651,
  164.6488,
  176.6236,
  167.0838,
  177.8864,
  162.6867,
  158.052,
  178.32,
  178.32,
  178.32,
  178.32,
  178.32,
  178.32 ;

 DZSOI =
  0.0175128188,
  0.0275789686,
  0.0454700328,
  0.0749674141,
  0.123600364,
  0.203782558,
  0.335980624,
  0.553938389,
  0.913290024,
  1.50576067,
  2.48257971,
  4.09308195,
  6.7483511,
  11.1261501,
  13.8511524 ;

 PCTSAND =
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000,
  20.000000;
															
 WATSAT =
  0.503309488,
  0.467856914,
  0.445469409,
  0.435835928,
  0.43314901,
  0.428174824,
  0.429554552,
  0.425283909,
  0.423480004,
  0.428519994,
  0.428519994,
  0.428519994,
  0.428519994,
  0.428519994,
  0.428519994 ;

 ZSOI =
  0.00710063521,
  0.0279249996,
  0.0622585751,
  0.118865065,
  0.2121934,
  0.3660658,
  0.619758487,
  1.03802705,
  1.72763526,
  2.8646071,
  4.73915672,
  7.82976627,
  12.9253206,
  21.3264694,
  35.1776199 ;

 lat = 38.8951988 ;

 levgrnd = 0.00710063521, 0.0279249996, 0.0622585751, 0.118865065, 0.2121934,
    0.3660658, 0.619758487, 1.03802705, 1.72763526, 2.8646071, 4.73915672,
    7.82976627, 12.9253206, 21.3264694, 35.1776199 ;

 lon = 239.367294 ;
}
